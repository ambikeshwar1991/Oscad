* EESchema Netlist Version 1.1 (Spice format) creation date: Thursday 01 August 2013 05:16:37 PM IST

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

*Sheet Name:/
U2  5 2 VPLOT8		
v2  4 0 DC		
U1  2 4 IPLOT		
D1  5 2 DIODE		
R1  1 5 100		
v1  1 0 SINE		

.end

* eeschema netlist version 1.1 (spice format) creation date: thursday 01 august 2013 05:16:37 pm ist

v2  4 0 dc 5
V_u1 2 4 0
d1  5 2 diode
r1  1 5 100
v1  1 0 sine(0 5 50 0 0)

.tran 10e-03 1e-01 0e-00
.plot v(5)-v(2) 
.plot i(V_u1)
.end

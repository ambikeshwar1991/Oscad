* eeschema netlist version 1.1 (spice format) creation date: monday 29 july 2013 01:04:39 pm ist
.include 1n4007.lib

* Plotting option vplot1
* Plotting option vplot
v1  in1 in2 sine(0 10 100 0 0)
c1  out gnd 1e-06
d4  gnd in2 1n4007
d2  in2 out 1n4007
d3  gnd in1 1n4007
d1  in1 out 1n4007
r1  out gnd 100000

.tran  100e-06 40e-03 0e-00
.plot v(out)
.plot v(in1)-v(in2)
.end

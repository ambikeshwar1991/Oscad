* EESchema Netlist Version 1.1 (Spice format) creation date: Monday 26 August 2013 12:32:59 PM IST

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

*Sheet Name:/
U1  8 vdbplot8_1		
v1  5 0 DC		
v2  2 0 AC		
R1  3 2 50		
R2  5 7 200k		
C1  3 7 40u		
R3  7 0 50k		
R6  8 0 1k		
C2  0 4 100u		
C3  8 6 40u		
R5  5 6 2k		
R4  4 0 1.5k		
Q1  4 7 6 NPN		

.end

* EESchema Netlist Version 1.1 (Spice format) creation date: Thursday 11 July 2013 05:13:06 PM IST

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

*Sheet Name:/
U1  N-000006 N-000007 N-000003 PORT		
Rout1  N-000003 N-000002 75		
Eout1  N-000002 GND N-000001 GND 1		
Cbw1  N-000001 GND 31.85e-9		
Rbw1  N-000001 N-000004 0.5e6		
Ein1  N-000004 GND N-000007 N-000006 100e3		
Rin1  N-000007 N-000006 2e6		

.end

* EESchema Netlist Version 1.1 (Spice format) creation date: Monday 29 July 2013 01:04:39 PM IST

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

*Sheet Name:/
U2  out VPLOT1		
U1  in1 in2 VPLOT		
V1  in1 in2 SINE		
C1  out GND 1e-06		
D4  GND in2 1n4007		
D2  in2 out 1n4007		
D3  GND in1 1n4007		
D1  in1 out 1n4007		
R1  out GND 100000		

.end

* eeschema netlist version 1.1 (spice format) creation date: monday 26 august 2013 12:32:59 pm ist
.include npn.lib

* Plotting option vdbplot8_1
v1  5 0 dc 10
v2  2 0 ac 1m
r1  3 2 50
r2  5 7 200k
c1  3 7 40u
r3  7 0 50k
r6  8 0 1k
c2  0 4 100u
c3  8 6 40u
r5  5 6 2k
r4  4 0 1.5k
q1 6 7 4 npn

.dc  v1 1e-00 4e-00 2e-00 v2 1e-00 5e-00 3e-00
.plot db(v(8)) 
.end
